library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.NUMERIC_STD.all;

entity tile_mem is
  port(
    tile_index : in unsigned(7 downto 0);
    tile_pixel_X : in unsigned(3 downto 0);
    tile_pixel_Y : in unsigned(3 downto 0);

    pixel_out : out unsigned(7 downto 0)
);
end tile_mem;

architecture Behavioral of tile_mem is
  type tMem_data is array (0 to 16383) of unsigned(7 downto 0);

  signal tMem : tMem_data :=
  (	--Black Tile
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",	
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",

	--Letter 0
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",	
    x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",
    x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",
    x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",
    x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",
    x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",
    x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",

	--Letter 1
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",

	--Letter 2
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",

	--Letter 3
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",

	--Letter 4
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",

	--Letter 5
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"FF",x"00",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"FF",x"FF",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",

	--Letter 6
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"FF",x"00",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"FF",x"FF",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",

	--Letter 7
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",

	--Letter 8
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",

	--Letter 9
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"FF",x"FF",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"FF",x"00",x"FF",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"FF",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",x"FF",x"FF",x"00",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",

        --Player Left
    x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",
    x"60",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"60",
    x"60",x"88",x"60",x"60",x"60",x"60",x"88",x"88",x"88",x"02",x"02",x"02",x"60",x"88",x"88",x"60",
    x"60",x"88",x"60",x"DF",x"DF",x"60",x"60",x"88",x"02",x"17",x"17",x"17",x"02",x"60",x"88",x"60",
    x"60",x"88",x"60",x"DF",x"DF",x"FF",x"FF",x"94",x"02",x"17",x"17",x"17",x"02",x"94",x"88",x"60",
    x"60",x"88",x"60",x"FF",x"FF",x"9F",x"FF",x"CC",x"02",x"17",x"17",x"17",x"02",x"CC",x"94",x"60",
    x"60",x"FF",x"FF",x"9F",x"93",x"9F",x"FF",x"CC",x"02",x"17",x"17",x"17",x"02",x"CC",x"94",x"60",
    x"FF",x"9F",x"93",x"9F",x"93",x"9F",x"FF",x"CC",x"CC",x"CC",x"CC",x"CC",x"CC",x"CC",x"94",x"60",
    x"60",x"FF",x"FF",x"9F",x"93",x"9F",x"94",x"94",x"94",x"94",x"94",x"94",x"94",x"94",x"88",x"60",
    x"60",x"88",x"88",x"FF",x"FF",x"94",x"40",x"40",x"40",x"AC",x"AC",x"40",x"40",x"40",x"94",x"60",
    x"60",x"88",x"88",x"88",x"88",x"94",x"40",x"AC",x"40",x"AC",x"AC",x"40",x"AC",x"40",x"94",x"60",
    x"60",x"88",x"88",x"88",x"88",x"94",x"40",x"40",x"40",x"AC",x"AC",x"40",x"40",x"40",x"94",x"60",
    x"60",x"88",x"88",x"88",x"88",x"60",x"94",x"94",x"94",x"94",x"94",x"94",x"94",x"94",x"88",x"60",
    x"60",x"88",x"88",x"88",x"88",x"60",x"60",x"60",x"60",x"88",x"88",x"88",x"88",x"88",x"88",x"60",
    x"60",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"60",
    x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",

        --Player Right
        x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",
        x"60",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"60",
        x"60",x"88",x"60",x"60",x"02",x"02",x"02",x"88",x"88",x"88",x"60",x"60",x"60",x"88",x"88",x"60",
        x"60",x"88",x"60",x"02",x"17",x"17",x"17",x"02",x"88",x"88",x"60",x"DF",x"60",x"60",x"88",x"60",
        x"60",x"88",x"94",x"02",x"17",x"17",x"17",x"02",x"94",x"FF",x"FF",x"DF",x"DF",x"60",x"88",x"60",
        x"60",x"94",x"CC",x"02",x"17",x"17",x"17",x"02",x"CC",x"FF",x"9F",x"FF",x"FF",x"60",x"88",x"60",
        x"60",x"94",x"CC",x"02",x"17",x"17",x"17",x"02",x"CC",x"FF",x"9F",x"93",x"9F",x"FF",x"FF",x"60",
        x"60",x"94",x"CC",x"CC",x"CC",x"CC",x"CC",x"CC",x"CC",x"FF",x"9F",x"93",x"9F",x"93",x"9F",x"FF",
        x"60",x"88",x"94",x"94",x"94",x"94",x"94",x"94",x"94",x"94",x"9F",x"93",x"9F",x"FF",x"FF",x"60",
        x"60",x"94",x"40",x"40",x"40",x"AC",x"AC",x"40",x"40",x"40",x"94",x"FF",x"FF",x"88",x"88",x"60",
        x"60",x"94",x"40",x"AC",x"40",x"AC",x"AC",x"40",x"AC",x"40",x"94",x"88",x"88",x"88",x"88",x"60",
        x"60",x"94",x"40",x"40",x"40",x"AC",x"AC",x"40",x"40",x"40",x"94",x"88",x"88",x"88",x"88",x"60",
        x"60",x"88",x"94",x"94",x"94",x"94",x"94",x"94",x"94",x"94",x"60",x"88",x"88",x"88",x"88",x"60",
        x"60",x"88",x"88",x"88",x"88",x"60",x"60",x"60",x"60",x"88",x"88",x"88",x"88",x"88",x"88",x"60",
        x"60",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"60",
        x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",

        --Player DOWN
    x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",
    x"60",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"60",
    x"60",x"88",x"60",x"94",x"94",x"60",x"88",x"02",x"02",x"02",x"60",x"60",x"94",x"94",x"88",x"60",
    x"60",x"88",x"60",x"94",x"94",x"CC",x"02",x"17",x"17",x"17",x"02",x"CC",x"94",x"94",x"88",x"60",
    x"60",x"88",x"60",x"94",x"94",x"CC",x"02",x"17",x"17",x"17",x"02",x"CC",x"94",x"94",x"88",x"60",
    x"60",x"88",x"60",x"94",x"94",x"CC",x"02",x"17",x"17",x"17",x"02",x"CC",x"94",x"94",x"88",x"60",
    x"60",x"88",x"88",x"94",x"94",x"CC",x"02",x"17",x"17",x"17",x"02",x"CC",x"94",x"94",x"88",x"60",
    x"60",x"88",x"88",x"94",x"94",x"CC",x"CC",x"CC",x"CC",x"CC",x"CC",x"CC",x"94",x"94",x"88",x"60",
    x"60",x"88",x"88",x"94",x"94",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"94",x"94",x"88",x"60",
    x"60",x"88",x"88",x"94",x"94",x"FF",x"9F",x"9F",x"9F",x"9F",x"9F",x"FF",x"94",x"94",x"88",x"60",
    x"60",x"88",x"88",x"94",x"94",x"60",x"FF",x"93",x"93",x"93",x"FF",x"88",x"94",x"94",x"88",x"60",
    x"60",x"88",x"88",x"88",x"88",x"60",x"FF",x"9F",x"9F",x"9F",x"FF",x"88",x"88",x"88",x"88",x"60",
    x"60",x"88",x"88",x"88",x"88",x"60",x"DF",x"FF",x"93",x"FF",x"88",x"88",x"88",x"88",x"88",x"60",
    x"60",x"88",x"88",x"88",x"88",x"60",x"60",x"FF",x"9F",x"FF",x"88",x"88",x"88",x"88",x"88",x"60",
    x"60",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"FF",x"88",x"88",x"88",x"88",x"88",x"88",x"60",
    x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",

        --Player UP
    x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",
    x"60",x"88",x"88",x"88",x"88",x"88",x"88",x"FF",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"60",
    x"60",x"88",x"60",x"60",x"60",x"60",x"FF",x"9F",x"FF",x"88",x"60",x"60",x"60",x"88",x"88",x"60",
    x"60",x"88",x"60",x"DF",x"DF",x"60",x"FF",x"93",x"FF",x"88",x"60",x"DF",x"60",x"60",x"88",x"60",
    x"60",x"88",x"60",x"DF",x"DF",x"FF",x"9F",x"9F",x"9F",x"FF",x"60",x"DF",x"DF",x"60",x"88",x"60",
    x"60",x"88",x"94",x"94",x"DF",x"FF",x"93",x"93",x"93",x"FF",x"60",x"94",x"94",x"60",x"88",x"60",
    x"60",x"88",x"94",x"94",x"FF",x"9F",x"02",x"02",x"02",x"9F",x"FF",x"94",x"94",x"60",x"88",x"60",
    x"60",x"88",x"94",x"94",x"FF",x"02",x"17",x"17",x"17",x"02",x"FF",x"94",x"94",x"60",x"88",x"60",
    x"60",x"88",x"94",x"94",x"CC",x"02",x"17",x"17",x"17",x"02",x"CC",x"94",x"94",x"60",x"88",x"60",
    x"60",x"88",x"94",x"94",x"CC",x"02",x"17",x"17",x"17",x"02",x"CC",x"94",x"94",x"88",x"88",x"60",
    x"60",x"88",x"94",x"94",x"CC",x"02",x"17",x"17",x"17",x"02",x"CC",x"94",x"94",x"88",x"88",x"60",
    x"60",x"88",x"94",x"94",x"CC",x"CC",x"CC",x"CC",x"CC",x"CC",x"CC",x"94",x"94",x"88",x"88",x"60",
    x"60",x"88",x"94",x"94",x"CC",x"CC",x"CC",x"CC",x"CC",x"CC",x"CC",x"94",x"94",x"88",x"88",x"60",
    x"60",x"88",x"94",x"94",x"88",x"60",x"60",x"60",x"60",x"88",x"88",x"94",x"94",x"88",x"88",x"60",
    x"60",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"60",
    x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",


        --BACKGROUND
    x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",
    x"60",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"60",
    x"60",x"88",x"60",x"60",x"60",x"60",x"88",x"88",x"88",x"88",x"60",x"60",x"60",x"88",x"88",x"60",
    x"60",x"88",x"60",x"DF",x"DF",x"60",x"60",x"88",x"88",x"88",x"60",x"DF",x"60",x"60",x"88",x"60",
    x"60",x"88",x"60",x"DF",x"DF",x"DF",x"60",x"88",x"88",x"88",x"60",x"DF",x"DF",x"60",x"88",x"60",
    x"60",x"88",x"60",x"60",x"DF",x"DF",x"60",x"88",x"88",x"88",x"60",x"60",x"DF",x"60",x"88",x"60",
    x"60",x"88",x"88",x"60",x"60",x"60",x"60",x"88",x"88",x"88",x"60",x"DF",x"DF",x"60",x"88",x"60",
    x"60",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"60",x"DF",x"DF",x"60",x"88",x"60",
    x"60",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"60",x"60",x"60",x"60",x"88",x"60",
    x"60",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"60",
    x"60",x"88",x"88",x"88",x"88",x"60",x"60",x"60",x"60",x"60",x"88",x"88",x"88",x"88",x"88",x"60",
    x"60",x"88",x"88",x"88",x"88",x"60",x"DF",x"DF",x"DF",x"60",x"88",x"88",x"88",x"88",x"88",x"60",
    x"60",x"88",x"88",x"88",x"88",x"60",x"DF",x"DF",x"60",x"60",x"88",x"88",x"88",x"88",x"88",x"60",
    x"60",x"88",x"88",x"88",x"88",x"60",x"60",x"60",x"60",x"88",x"88",x"88",x"88",x"88",x"88",x"60",
    x"60",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"88",x"60",
    x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",

        --THE ROCK
    x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",
    x"60",x"60",x"60",x"60",x"77",x"77",x"77",x"77",x"77",x"77",x"77",x"77",x"60",x"60",x"60",x"60",
    x"60",x"60",x"77",x"77",x"77",x"B6",x"B6",x"B6",x"B6",x"B6",x"B6",x"77",x"77",x"77",x"60",x"60",
    x"60",x"60",x"77",x"B6",x"B6",x"B6",x"B6",x"B6",x"B6",x"B6",x"B6",x"B6",x"B6",x"77",x"60",x"60",
    x"60",x"77",x"77",x"B6",x"B6",x"B6",x"B6",x"B6",x"B6",x"B6",x"B6",x"B6",x"B6",x"77",x"77",x"60",
    x"60",x"77",x"B6",x"B6",x"B6",x"B6",x"B6",x"B6",x"B6",x"B6",x"B6",x"B6",x"B6",x"B6",x"77",x"60",
    x"60",x"77",x"B6",x"B6",x"B6",x"B6",x"B6",x"B6",x"B6",x"B6",x"B6",x"B6",x"B6",x"B6",x"77",x"60",
    x"60",x"77",x"B6",x"B6",x"B6",x"B6",x"B6",x"B6",x"B6",x"B6",x"B6",x"B6",x"B6",x"B6",x"77",x"60",
    x"60",x"77",x"B6",x"B6",x"B6",x"B6",x"B6",x"B6",x"B6",x"B6",x"B6",x"B6",x"B6",x"B6",x"77",x"60",
    x"60",x"77",x"B6",x"B6",x"B6",x"B6",x"B6",x"B6",x"B6",x"B6",x"B6",x"B6",x"B6",x"B6",x"77",x"60",
    x"60",x"77",x"B6",x"B6",x"B6",x"B6",x"B6",x"B6",x"B6",x"B6",x"B6",x"B6",x"B6",x"B6",x"77",x"60",
    x"60",x"77",x"77",x"B6",x"B6",x"B6",x"B6",x"B6",x"B6",x"B6",x"B6",x"B6",x"B6",x"77",x"77",x"60",
    x"60",x"60",x"77",x"B6",x"B6",x"B6",x"B6",x"B6",x"B6",x"B6",x"B6",x"B6",x"B6",x"77",x"60",x"60",
    x"60",x"60",x"77",x"77",x"77",x"B6",x"B6",x"B6",x"B6",x"B6",x"B6",x"77",x"77",x"77",x"60",x"60",
    x"60",x"60",x"60",x"60",x"77",x"77",x"77",x"77",x"77",x"77",x"77",x"77",x"60",x"60",x"60",x"60",
    x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",

        --THE ROCK OF SILVER
    x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",
    x"60",x"60",x"60",x"60",x"77",x"77",x"77",x"77",x"77",x"77",x"77",x"77",x"60",x"60",x"60",x"60",
    x"60",x"60",x"77",x"77",x"77",x"B6",x"B6",x"B6",x"B6",x"B6",x"B6",x"77",x"77",x"77",x"60",x"60",
    x"60",x"60",x"77",x"B6",x"B6",x"B6",x"B6",x"B6",x"B6",x"B6",x"B6",x"B6",x"B6",x"77",x"60",x"60",
    x"60",x"77",x"77",x"B6",x"B6",x"7B",x"B6",x"B6",x"B6",x"B6",x"B6",x"B6",x"B6",x"77",x"77",x"60",
    x"60",x"77",x"B6",x"B6",x"B6",x"7B",x"B6",x"B6",x"B6",x"7B",x"7B",x"B6",x"B6",x"B6",x"77",x"60",
    x"60",x"77",x"B6",x"B6",x"7B",x"7B",x"B6",x"B6",x"B6",x"B6",x"7B",x"7B",x"7B",x"B6",x"77",x"60",
    x"60",x"77",x"B6",x"B6",x"7B",x"B6",x"B6",x"B6",x"B6",x"B6",x"B6",x"B6",x"7B",x"B6",x"77",x"60",
    x"60",x"77",x"B6",x"B6",x"B6",x"B6",x"B6",x"B6",x"B6",x"B6",x"B6",x"B6",x"7B",x"B6",x"77",x"60",
    x"60",x"77",x"B6",x"B6",x"B6",x"B6",x"7B",x"7B",x"7B",x"B6",x"B6",x"B6",x"B6",x"B6",x"77",x"60",
    x"60",x"77",x"B6",x"B6",x"B6",x"7B",x"7B",x"B6",x"7B",x"7B",x"7B",x"B6",x"B6",x"B6",x"77",x"60",
    x"60",x"77",x"77",x"B6",x"B6",x"B6",x"B6",x"B6",x"B6",x"B6",x"B6",x"B6",x"B6",x"77",x"77",x"60",
    x"60",x"60",x"77",x"B6",x"B6",x"B6",x"B6",x"B6",x"B6",x"B6",x"B6",x"B6",x"B6",x"77",x"60",x"60",
    x"60",x"60",x"77",x"77",x"77",x"B6",x"B6",x"B6",x"B6",x"B6",x"B6",x"77",x"77",x"77",x"60",x"60",
    x"60",x"60",x"60",x"60",x"77",x"77",x"77",x"77",x"77",x"77",x"77",x"77",x"60",x"60",x"60",x"60",
    x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",

       --THE ROCK OF GOLD
    x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",
    x"60",x"60",x"60",x"60",x"77",x"77",x"77",x"77",x"77",x"77",x"77",x"77",x"60",x"60",x"60",x"60",
    x"60",x"60",x"77",x"77",x"77",x"B6",x"B6",x"B6",x"B6",x"B6",x"B6",x"77",x"77",x"77",x"60",x"60",
    x"60",x"60",x"77",x"B6",x"B6",x"B6",x"B6",x"B6",x"B6",x"B6",x"B6",x"B6",x"B6",x"77",x"60",x"60",
    x"60",x"77",x"77",x"B6",x"B6",x"DD",x"B6",x"B6",x"B6",x"B6",x"B6",x"B6",x"B6",x"77",x"77",x"60",
    x"60",x"77",x"B6",x"B6",x"B6",x"DD",x"B6",x"B6",x"B6",x"DD",x"DD",x"B6",x"B6",x"B6",x"77",x"60",
    x"60",x"77",x"B6",x"B6",x"DD",x"DD",x"B6",x"B6",x"B6",x"B6",x"DD",x"DD",x"DD",x"B6",x"77",x"60",
    x"60",x"77",x"B6",x"B6",x"DD",x"B6",x"B6",x"B6",x"B6",x"B6",x"B6",x"B6",x"DD",x"B6",x"77",x"60",
    x"60",x"77",x"B6",x"B6",x"B6",x"B6",x"B6",x"B6",x"B6",x"B6",x"B6",x"B6",x"DD",x"B6",x"77",x"60",
    x"60",x"77",x"B6",x"B6",x"B6",x"B6",x"DD",x"DD",x"DD",x"B6",x"B6",x"B6",x"B6",x"B6",x"77",x"60",
    x"60",x"77",x"B6",x"B6",x"B6",x"DD",x"DD",x"B6",x"DD",x"DD",x"DD",x"B6",x"B6",x"B6",x"77",x"60",
    x"60",x"77",x"77",x"B6",x"B6",x"B6",x"B6",x"B6",x"B6",x"B6",x"B6",x"B6",x"B6",x"77",x"77",x"60",
    x"60",x"60",x"77",x"B6",x"B6",x"B6",x"B6",x"B6",x"B6",x"B6",x"B6",x"B6",x"B6",x"77",x"60",x"60",
    x"60",x"60",x"77",x"77",x"77",x"B6",x"B6",x"B6",x"B6",x"B6",x"B6",x"77",x"77",x"77",x"60",x"60",
    x"60",x"60",x"60",x"60",x"77",x"77",x"77",x"77",x"77",x"77",x"77",x"77",x"60",x"60",x"60",x"60",
    x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",

      --THE ROCK OF greed
    x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",
    x"60",x"60",x"60",x"60",x"77",x"77",x"77",x"77",x"77",x"77",x"77",x"77",x"60",x"60",x"60",x"60",
    x"60",x"60",x"77",x"77",x"77",x"B6",x"B6",x"B6",x"B6",x"B6",x"B6",x"77",x"77",x"77",x"60",x"60",
    x"60",x"60",x"77",x"B6",x"B6",x"B6",x"B6",x"B6",x"B6",x"B6",x"B6",x"B6",x"B6",x"77",x"60",x"60",
    x"60",x"77",x"77",x"B6",x"B6",x"B6",x"B6",x"B6",x"B6",x"E4",x"E4",x"B6",x"B6",x"77",x"77",x"60",
    x"60",x"77",x"B6",x"B6",x"E4",x"B6",x"B6",x"B6",x"E4",x"C0",x"C0",x"E4",x"B6",x"B6",x"77",x"60",
    x"60",x"77",x"B6",x"E4",x"C0",x"E4",x"B6",x"B6",x"E4",x"C0",x"C0",x"E4",x"B6",x"B6",x"77",x"60",
    x"60",x"77",x"B6",x"E4",x"C0",x"E4",x"B6",x"B6",x"E4",x"C0",x"C0",x"E4",x"B6",x"B6",x"77",x"60",
    x"60",x"77",x"B6",x"B6",x"E4",x"B6",x"B6",x"B6",x"B6",x"E4",x"E4",x"B6",x"B6",x"B6",x"77",x"60",
    x"60",x"77",x"B6",x"B6",x"B6",x"B6",x"B6",x"B6",x"B6",x"B6",x"B6",x"B6",x"B6",x"B6",x"77",x"60",
    x"60",x"77",x"B6",x"B6",x"B6",x"B6",x"E4",x"E4",x"E4",x"B6",x"B6",x"B6",x"B6",x"B6",x"77",x"60",
    x"60",x"77",x"77",x"B6",x"B6",x"E4",x"C0",x"C0",x"C0",x"E4",x"B6",x"B6",x"B6",x"77",x"77",x"60",
    x"60",x"60",x"77",x"B6",x"B6",x"B6",x"E4",x"E4",x"E4",x"B6",x"B6",x"B6",x"B6",x"77",x"60",x"60",
    x"60",x"60",x"77",x"77",x"77",x"B6",x"B6",x"B6",x"B6",x"B6",x"B6",x"77",x"77",x"77",x"60",x"60",
    x"60",x"60",x"60",x"60",x"77",x"77",x"77",x"77",x"77",x"77",x"77",x"77",x"60",x"60",x"60",x"60",
    x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",

    --Drill Icon
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"00",x"00",x"00",
    x"00",x"00",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"00",x"00",
    x"00",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"00",  
    x"00",x"EC",x"EC",x"00",x"00",x"00",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"00",
    x"00",x"EC",x"EC",x"00",x"9F",x"9F",x"00",x"00",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"00",
    x"00",x"EC",x"EC",x"00",x"9F",x"9F",x"93",x"93",x"00",x"00",x"EC",x"EC",x"EC",x"EC",x"EC",x"00",
    x"00",x"EC",x"EC",x"00",x"9F",x"9F",x"93",x"93",x"9F",x"9F",x"00",x"00",x"EC",x"EC",x"EC",x"00",
    x"00",x"EC",x"EC",x"00",x"9F",x"93",x"93",x"9F",x"9F",x"93",x"93",x"9F",x"00",x"00",x"EC",x"00",
    x"00",x"EC",x"EC",x"00",x"9F",x"93",x"93",x"9F",x"9F",x"93",x"00",x"00",x"EC",x"EC",x"EC",x"00",
    x"00",x"EC",x"EC",x"00",x"9F",x"93",x"93",x"9F",x"00",x"00",x"EC",x"EC",x"EC",x"EC",x"EC",x"00",
    x"00",x"EC",x"EC",x"00",x"93",x"93",x"00",x"00",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"00",  
    x"00",x"EC",x"EC",x"00",x"00",x"00",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"00",
    x"00",x"00",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"00",x"00",
    x"00",x"00",x"00",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"EC",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",

        --Peng Icon          
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"00",x"00",x"00",
    x"00",x"00",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"00",x"00",
    x"00",x"FC",x"FC",x"FC",x"FC",x"FC",x"1C",x"1C",x"1C",x"1C",x"1C",x"FC",x"FC",x"FC",x"FC",x"00",
    x"00",x"FC",x"FC",x"FC",x"FC",x"FC",x"1C",x"1C",x"FC",x"FC",x"FC",x"1C",x"FC",x"FC",x"FC",x"00",
    x"00",x"FC",x"FC",x"FC",x"FC",x"FC",x"1C",x"1C",x"FC",x"FC",x"FC",x"1C",x"FC",x"FC",x"FC",x"00",
    x"00",x"FC",x"FC",x"FC",x"FC",x"FC",x"1C",x"1C",x"FC",x"FC",x"FC",x"1C",x"FC",x"FC",x"FC",x"00",
    x"00",x"FC",x"FC",x"FC",x"FC",x"FC",x"1C",x"1C",x"FC",x"FC",x"FC",x"1C",x"FC",x"FC",x"FC",x"00",
    x"00",x"FC",x"FC",x"FC",x"FC",x"FC",x"1C",x"1C",x"1C",x"1C",x"1C",x"FC",x"FC",x"FC",x"FC",x"00",
    x"00",x"FC",x"FC",x"FC",x"FC",x"FC",x"1C",x"1C",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"00",
    x"00",x"FC",x"FC",x"FC",x"FC",x"1C",x"1C",x"1C",x"1C",x"1C",x"FC",x"FC",x"FC",x"FC",x"FC",x"00",
    x"00",x"FC",x"FC",x"FC",x"FC",x"FC",x"1C",x"1C",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"00",
    x"00",x"FC",x"FC",x"FC",x"FC",x"1C",x"1C",x"1C",x"1C",x"1C",x"FC",x"FC",x"FC",x"FC",x"FC",x"00",
    x"00",x"00",x"FC",x"FC",x"FC",x"FC",x"1C",x"1C",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"00",x"00",
    x"00",x"00",x"00",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",    

        --Icon template      
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
    x"00",x"00",x"00",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"00",x"00",x"00",
    x"00",x"00",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"00",x"00",
    x"00",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"00",
    x"00",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"00",
    x"00",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"00",
    x"00",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"00",
    x"00",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"00",
    x"00",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"00",
    x"00",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"00",
    x"00",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"00",
    x"00",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"00",
    x"00",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"00",
    x"00",x"00",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"00",x"00",
    x"00",x"00",x"00",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"FC",x"00",x"00",x"00",
    x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",
        
x"30",x"30",x"30",x"30",x"31",x"31",x"31",x"31",x"32",x"32",x"32",x"32",x"33",x"33",x"33",x"33",
x"30",x"30",x"30",x"30",x"31",x"31",x"31",x"31",x"32",x"32",x"32",x"32",x"33",x"33",x"33",x"33",
x"30",x"30",x"30",x"30",x"31",x"31",x"31",x"31",x"32",x"32",x"32",x"32",x"33",x"33",x"33",x"33",
x"30",x"30",x"30",x"30",x"31",x"31",x"31",x"31",x"32",x"32",x"32",x"32",x"33",x"33",x"33",x"33",
x"34",x"34",x"34",x"34",x"35",x"35",x"35",x"35",x"36",x"36",x"36",x"36",x"37",x"37",x"37",x"37",
x"34",x"34",x"34",x"34",x"35",x"35",x"35",x"35",x"36",x"36",x"36",x"36",x"37",x"37",x"37",x"37",
x"34",x"34",x"34",x"34",x"35",x"35",x"35",x"35",x"36",x"36",x"36",x"36",x"37",x"37",x"37",x"37",
x"34",x"34",x"34",x"34",x"35",x"35",x"35",x"35",x"36",x"36",x"36",x"36",x"37",x"37",x"37",x"37",
x"38",x"38",x"38",x"38",x"39",x"39",x"39",x"39",x"3A",x"3A",x"3A",x"3A",x"3B",x"3B",x"3B",x"3B",
x"38",x"38",x"38",x"38",x"39",x"39",x"39",x"39",x"3A",x"3A",x"3A",x"3A",x"3B",x"3B",x"3B",x"3B",
x"38",x"38",x"38",x"38",x"39",x"39",x"39",x"39",x"3A",x"3A",x"3A",x"3A",x"3B",x"3B",x"3B",x"3B",
x"38",x"38",x"38",x"38",x"39",x"39",x"39",x"39",x"3A",x"3A",x"3A",x"3A",x"3B",x"3B",x"3B",x"3B",
x"3C",x"3C",x"3C",x"3C",x"3D",x"3D",x"3D",x"3D",x"3E",x"3E",x"3E",x"3E",x"3F",x"3F",x"3F",x"3F",
x"3C",x"3C",x"3C",x"3C",x"3D",x"3D",x"3D",x"3D",x"3E",x"3E",x"3E",x"3E",x"3F",x"3F",x"3F",x"3F",
x"3C",x"3C",x"3C",x"3C",x"3D",x"3D",x"3D",x"3D",x"3E",x"3E",x"3E",x"3E",x"3F",x"3F",x"3F",x"3F",
x"3C",x"3C",x"3C",x"3C",x"3D",x"3D",x"3D",x"3D",x"3E",x"3E",x"3E",x"3E",x"3F",x"3F",x"3F",x"3F",


x"40",x"40",x"40",x"40",x"41",x"41",x"41",x"41",x"42",x"42",x"42",x"42",x"77",x"77",x"77",x"77",
x"40",x"40",x"40",x"40",x"41",x"41",x"41",x"41",x"42",x"42",x"42",x"42",x"77",x"77",x"77",x"77",
x"40",x"40",x"40",x"40",x"41",x"41",x"41",x"41",x"42",x"42",x"42",x"42",x"77",x"77",x"77",x"77",
x"40",x"40",x"40",x"40",x"41",x"41",x"41",x"41",x"42",x"42",x"42",x"42",x"77",x"77",x"77",x"77",
x"44",x"44",x"44",x"44",x"45",x"45",x"45",x"45",x"46",x"46",x"46",x"46",x"47",x"47",x"47",x"47",
x"44",x"44",x"44",x"44",x"45",x"45",x"45",x"45",x"46",x"46",x"46",x"46",x"47",x"47",x"47",x"47",
x"44",x"44",x"44",x"44",x"45",x"45",x"45",x"45",x"46",x"46",x"46",x"46",x"47",x"47",x"47",x"47",
x"44",x"44",x"44",x"44",x"45",x"45",x"45",x"45",x"46",x"46",x"46",x"46",x"47",x"47",x"47",x"47",
x"48",x"48",x"48",x"48",x"49",x"49",x"49",x"49",x"4A",x"4A",x"4A",x"4A",x"4B",x"4B",x"4B",x"4B",
x"48",x"48",x"48",x"48",x"49",x"49",x"49",x"49",x"4A",x"4A",x"4A",x"4A",x"4B",x"4B",x"4B",x"4B",
x"48",x"48",x"48",x"48",x"49",x"49",x"49",x"49",x"4A",x"4A",x"4A",x"4A",x"4B",x"4B",x"4B",x"4B",
x"48",x"48",x"48",x"48",x"49",x"49",x"49",x"49",x"4A",x"4A",x"4A",x"4A",x"4B",x"4B",x"4B",x"4B",
x"4C",x"4C",x"4C",x"4C",x"4D",x"4D",x"4D",x"4D",x"4E",x"4E",x"4E",x"4E",x"4F",x"4F",x"4F",x"4F",
x"4C",x"4C",x"4C",x"4C",x"4D",x"4D",x"4D",x"4D",x"4E",x"4E",x"4E",x"4E",x"4F",x"4F",x"4F",x"4F",
x"4C",x"4C",x"4C",x"4C",x"4D",x"4D",x"4D",x"4D",x"4E",x"4E",x"4E",x"4E",x"4F",x"4F",x"4F",x"4F",
x"4C",x"4C",x"4C",x"4C",x"4D",x"4D",x"4D",x"4D",x"4E",x"4E",x"4E",x"4E",x"4F",x"4F",x"4F",x"4F",


x"50",x"50",x"50",x"50",x"51",x"51",x"51",x"51",x"52",x"52",x"52",x"52",x"53",x"53",x"53",x"53",
x"50",x"50",x"50",x"50",x"51",x"51",x"51",x"51",x"52",x"52",x"52",x"52",x"53",x"53",x"53",x"53",
x"50",x"50",x"50",x"50",x"51",x"51",x"51",x"51",x"52",x"52",x"52",x"52",x"53",x"53",x"53",x"53",
x"50",x"50",x"50",x"50",x"51",x"51",x"51",x"51",x"52",x"52",x"52",x"52",x"53",x"53",x"53",x"53",
x"54",x"54",x"54",x"54",x"55",x"55",x"55",x"55",x"56",x"56",x"56",x"56",x"57",x"57",x"57",x"57",
x"54",x"54",x"54",x"54",x"55",x"55",x"55",x"55",x"56",x"56",x"56",x"56",x"57",x"57",x"57",x"57",
x"54",x"54",x"54",x"54",x"55",x"55",x"55",x"55",x"56",x"56",x"56",x"56",x"57",x"57",x"57",x"57",
x"54",x"54",x"54",x"54",x"55",x"55",x"55",x"55",x"56",x"56",x"56",x"56",x"57",x"57",x"57",x"57",
x"58",x"58",x"58",x"58",x"59",x"59",x"59",x"59",x"5A",x"5A",x"5A",x"5A",x"5B",x"5B",x"5B",x"5B",
x"58",x"58",x"58",x"58",x"59",x"59",x"59",x"59",x"5A",x"5A",x"5A",x"5A",x"5B",x"5B",x"5B",x"5B",
x"58",x"58",x"58",x"58",x"59",x"59",x"59",x"59",x"5A",x"5A",x"5A",x"5A",x"5B",x"5B",x"5B",x"5B",
x"58",x"58",x"58",x"58",x"59",x"59",x"59",x"59",x"5A",x"5A",x"5A",x"5A",x"5B",x"5B",x"5B",x"5B",
x"5C",x"5C",x"5C",x"5C",x"5D",x"5D",x"5D",x"5D",x"5E",x"5E",x"5E",x"5E",x"5F",x"5F",x"5F",x"5F",
x"5C",x"5C",x"5C",x"5C",x"5D",x"5D",x"5D",x"5D",x"5E",x"5E",x"5E",x"5E",x"5F",x"5F",x"5F",x"5F",
x"5C",x"5C",x"5C",x"5C",x"5D",x"5D",x"5D",x"5D",x"5E",x"5E",x"5E",x"5E",x"5F",x"5F",x"5F",x"5F",
x"5C",x"5C",x"5C",x"5C",x"5D",x"5D",x"5D",x"5D",x"5E",x"5E",x"5E",x"5E",x"5F",x"5F",x"5F",x"5F",


x"60",x"60",x"60",x"60",x"61",x"61",x"61",x"61",x"62",x"62",x"62",x"62",x"63",x"63",x"63",x"63",
x"60",x"60",x"60",x"60",x"61",x"61",x"61",x"61",x"62",x"62",x"62",x"62",x"63",x"63",x"63",x"63",
x"60",x"60",x"60",x"60",x"61",x"61",x"61",x"61",x"62",x"62",x"62",x"62",x"63",x"63",x"63",x"63",
x"60",x"60",x"60",x"60",x"61",x"61",x"61",x"61",x"62",x"62",x"62",x"62",x"63",x"63",x"63",x"63",
x"64",x"64",x"64",x"64",x"65",x"65",x"65",x"65",x"66",x"66",x"66",x"66",x"67",x"67",x"67",x"67",
x"64",x"64",x"64",x"64",x"65",x"65",x"65",x"65",x"66",x"66",x"66",x"66",x"67",x"67",x"67",x"67",
x"64",x"64",x"64",x"64",x"65",x"65",x"65",x"65",x"66",x"66",x"66",x"66",x"67",x"67",x"67",x"67",
x"64",x"64",x"64",x"64",x"65",x"65",x"65",x"65",x"66",x"66",x"66",x"66",x"67",x"67",x"67",x"67",
x"68",x"68",x"68",x"68",x"69",x"69",x"69",x"69",x"6A",x"6A",x"6A",x"6A",x"6B",x"6B",x"6B",x"6B",
x"68",x"68",x"68",x"68",x"69",x"69",x"69",x"69",x"6A",x"6A",x"6A",x"6A",x"6B",x"6B",x"6B",x"6B",
x"68",x"68",x"68",x"68",x"69",x"69",x"69",x"69",x"6A",x"6A",x"6A",x"6A",x"6B",x"6B",x"6B",x"6B",
x"68",x"68",x"68",x"68",x"69",x"69",x"69",x"69",x"6A",x"6A",x"6A",x"6A",x"6B",x"6B",x"6B",x"6B",
x"6C",x"6C",x"6C",x"6C",x"6D",x"6D",x"6D",x"6D",x"6E",x"6E",x"6E",x"6E",x"6F",x"6F",x"6F",x"6F",
x"6C",x"6C",x"6C",x"6C",x"6D",x"6D",x"6D",x"6D",x"6E",x"6E",x"6E",x"6E",x"6F",x"6F",x"6F",x"6F",
x"6C",x"6C",x"6C",x"6C",x"6D",x"6D",x"6D",x"6D",x"6E",x"6E",x"6E",x"6E",x"6F",x"6F",x"6F",x"6F",
x"6C",x"6C",x"6C",x"6C",x"6D",x"6D",x"6D",x"6D",x"6E",x"6E",x"6E",x"6E",x"6F",x"6F",x"6F",x"6F",


x"70",x"70",x"70",x"70",x"71",x"71",x"71",x"71",x"72",x"72",x"72",x"72",x"DF",x"DF",x"DF",x"DF",
x"70",x"70",x"70",x"70",x"71",x"71",x"71",x"71",x"72",x"72",x"72",x"72",x"DF",x"DF",x"DF",x"DF",
x"70",x"70",x"70",x"70",x"71",x"71",x"71",x"71",x"72",x"72",x"72",x"72",x"DF",x"DF",x"DF",x"DF",
x"70",x"70",x"70",x"70",x"71",x"71",x"71",x"71",x"72",x"72",x"72",x"72",x"DF",x"DF",x"DF",x"DF",
x"74",x"74",x"74",x"74",x"75",x"75",x"75",x"75",x"76",x"76",x"76",x"76",x"DF",x"DF",x"DF",x"DF",
x"74",x"74",x"74",x"74",x"75",x"75",x"75",x"75",x"76",x"76",x"76",x"76",x"DF",x"DF",x"DF",x"DF",
x"74",x"74",x"74",x"74",x"75",x"75",x"75",x"75",x"76",x"76",x"76",x"76",x"DF",x"DF",x"DF",x"DF",
x"74",x"74",x"74",x"74",x"75",x"75",x"75",x"75",x"76",x"76",x"76",x"76",x"DF",x"DF",x"DF",x"DF",
x"78",x"78",x"78",x"78",x"79",x"79",x"79",x"79",x"7A",x"7A",x"7A",x"7A",x"7B",x"7B",x"7B",x"7B",
x"78",x"78",x"78",x"78",x"79",x"79",x"79",x"79",x"7A",x"7A",x"7A",x"7A",x"7B",x"7B",x"7B",x"7B",
x"78",x"78",x"78",x"78",x"79",x"79",x"79",x"79",x"7A",x"7A",x"7A",x"7A",x"7B",x"7B",x"7B",x"7B",
x"78",x"78",x"78",x"78",x"79",x"79",x"79",x"79",x"7A",x"7A",x"7A",x"7A",x"7B",x"7B",x"7B",x"7B",
x"7C",x"7C",x"7C",x"7C",x"7D",x"7D",x"7D",x"7D",x"7E",x"7E",x"7E",x"7E",x"7F",x"7F",x"7F",x"7F",
x"7C",x"7C",x"7C",x"7C",x"7D",x"7D",x"7D",x"7D",x"7E",x"7E",x"7E",x"7E",x"7F",x"7F",x"7F",x"7F",
x"7C",x"7C",x"7C",x"7C",x"7D",x"7D",x"7D",x"7D",x"7E",x"7E",x"7E",x"7E",x"7F",x"7F",x"7F",x"7F",
x"7C",x"7C",x"7C",x"7C",x"7D",x"7D",x"7D",x"7D",x"7E",x"7E",x"7E",x"7E",x"7F",x"7F",x"7F",x"7F",


x"80",x"80",x"80",x"80",x"81",x"81",x"81",x"81",x"82",x"82",x"82",x"82",x"83",x"83",x"83",x"83",
x"80",x"80",x"80",x"80",x"81",x"81",x"81",x"81",x"82",x"82",x"82",x"82",x"83",x"83",x"83",x"83",
x"80",x"80",x"80",x"80",x"81",x"81",x"81",x"81",x"82",x"82",x"82",x"82",x"83",x"83",x"83",x"83",
x"80",x"80",x"80",x"80",x"81",x"81",x"81",x"81",x"82",x"82",x"82",x"82",x"83",x"83",x"83",x"83",
x"84",x"84",x"84",x"84",x"85",x"85",x"85",x"85",x"86",x"86",x"86",x"86",x"87",x"87",x"87",x"87",
x"84",x"84",x"84",x"84",x"85",x"85",x"85",x"85",x"86",x"86",x"86",x"86",x"87",x"87",x"87",x"87",
x"84",x"84",x"84",x"84",x"85",x"85",x"85",x"85",x"86",x"86",x"86",x"86",x"87",x"87",x"87",x"87",
x"84",x"84",x"84",x"84",x"85",x"85",x"85",x"85",x"86",x"86",x"86",x"86",x"87",x"87",x"87",x"87",
x"88",x"88",x"88",x"88",x"89",x"89",x"89",x"89",x"8A",x"8A",x"8A",x"8A",x"8B",x"8B",x"8B",x"8B",
x"88",x"88",x"88",x"88",x"89",x"89",x"89",x"89",x"8A",x"8A",x"8A",x"8A",x"8B",x"8B",x"8B",x"8B",
x"88",x"88",x"88",x"88",x"89",x"89",x"89",x"89",x"8A",x"8A",x"8A",x"8A",x"8B",x"8B",x"8B",x"8B",
x"88",x"88",x"88",x"88",x"89",x"89",x"89",x"89",x"8A",x"8A",x"8A",x"8A",x"8B",x"8B",x"8B",x"8B",
x"8C",x"8C",x"8C",x"8C",x"8D",x"8D",x"8D",x"8D",x"8E",x"8E",x"8E",x"8E",x"8F",x"8F",x"8F",x"8F",
x"8C",x"8C",x"8C",x"8C",x"8D",x"8D",x"8D",x"8D",x"8E",x"8E",x"8E",x"8E",x"8F",x"8F",x"8F",x"8F",
x"8C",x"8C",x"8C",x"8C",x"8D",x"8D",x"8D",x"8D",x"8E",x"8E",x"8E",x"8E",x"8F",x"8F",x"8F",x"8F",
x"8C",x"8C",x"8C",x"8C",x"8D",x"8D",x"8D",x"8D",x"8E",x"8E",x"8E",x"8E",x"8F",x"8F",x"8F",x"8F",

--Cracked Rocks (HEX adress = ??)
    x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",
    x"60",x"60",x"60",x"60",x"77",x"77",x"00",x"77",x"77",x"77",x"77",x"77",x"60",x"60",x"60",x"60",
    x"60",x"60",x"77",x"00",x"00",x"B6",x"00",x"B6",x"B6",x"B6",x"B6",x"00",x"77",x"77",x"60",x"60",
    x"60",x"60",x"77",x"B6",x"B6",x"00",x"00",x"B6",x"B6",x"00",x"00",x"B6",x"B6",x"77",x"60",x"60",
    x"60",x"77",x"00",x"B6",x"00",x"B6",x"B6",x"00",x"00",x"B6",x"B6",x"B6",x"B6",x"77",x"77",x"60",
    x"60",x"77",x"B6",x"00",x"B6",x"B6",x"B6",x"00",x"B6",x"B6",x"B6",x"B6",x"B6",x"00",x"00",x"60",
    x"60",x"77",x"B6",x"B6",x"B6",x"B6",x"00",x"B6",x"B6",x"B6",x"B6",x"B6",x"00",x"B6",x"77",x"60",
    x"60",x"77",x"B6",x"B6",x"B6",x"B6",x"00",x"B6",x"B6",x"B6",x"B6",x"00",x"00",x"B6",x"77",x"60",
    x"60",x"77",x"B6",x"B6",x"B6",x"B6",x"00",x"B6",x"B6",x"B6",x"B6",x"B6",x"B6",x"00",x"77",x"60",
    x"60",x"00",x"B6",x"B6",x"B6",x"00",x"B6",x"00",x"00",x"B6",x"B6",x"B6",x"B6",x"00",x"77",x"60",
    x"60",x"77",x"00",x"B6",x"B6",x"00",x"B6",x"B6",x"B6",x"00",x"B6",x"B6",x"00",x"B6",x"77",x"60",
    x"60",x"77",x"00",x"B6",x"00",x"B6",x"B6",x"B6",x"B6",x"B6",x"00",x"B6",x"00",x"77",x"77",x"60",
    x"60",x"60",x"77",x"00",x"B6",x"B6",x"B6",x"B6",x"B6",x"B6",x"B6",x"00",x"B6",x"00",x"60",x"60",
    x"60",x"60",x"77",x"00",x"77",x"B6",x"B6",x"00",x"B6",x"B6",x"B6",x"00",x"77",x"77",x"60",x"60",
    x"60",x"60",x"60",x"60",x"77",x"77",x"77",x"00",x"77",x"77",x"00",x"77",x"60",x"60",x"60",x"60",
    x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",

        --THE CRACKED ROCK OF SILVER
    x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",
    x"60",x"60",x"60",x"60",x"77",x"77",x"00",x"77",x"77",x"77",x"77",x"77",x"60",x"60",x"60",x"60",
    x"60",x"60",x"77",x"00",x"00",x"B6",x"00",x"B6",x"B6",x"B6",x"B6",x"00",x"77",x"77",x"60",x"60",
    x"60",x"60",x"77",x"B6",x"B6",x"00",x"00",x"B6",x"B6",x"00",x"00",x"B6",x"B6",x"77",x"60",x"60",
    x"60",x"77",x"00",x"B6",x"00",x"7B",x"B6",x"00",x"00",x"B6",x"B6",x"B6",x"B6",x"77",x"77",x"60",
    x"60",x"77",x"B6",x"00",x"B6",x"7B",x"B6",x"00",x"B6",x"7B",x"7B",x"B6",x"B6",x"00",x"00",x"60",
    x"60",x"77",x"B6",x"B6",x"7B",x"7B",x"00",x"B6",x"B6",x"B6",x"7B",x"7B",x"00",x"B6",x"77",x"60",
    x"60",x"77",x"B6",x"B6",x"7B",x"B6",x"00",x"B6",x"B6",x"B6",x"B6",x"00",x"00",x"B6",x"77",x"60",
    x"60",x"77",x"B6",x"B6",x"B6",x"B6",x"00",x"B6",x"B6",x"B6",x"B6",x"B6",x"7B",x"00",x"77",x"60",
    x"60",x"77",x"B6",x"B6",x"B6",x"00",x"7B",x"00",x"00",x"B6",x"B6",x"B6",x"B6",x"00",x"77",x"60",
    x"60",x"00",x"00",x"B6",x"B6",x"00",x"7B",x"B6",x"7B",x"00",x"7B",x"B6",x"00",x"B6",x"77",x"60",
    x"60",x"77",x"00",x"B6",x"00",x"B6",x"B6",x"B6",x"B6",x"B6",x"00",x"B6",x"00",x"77",x"77",x"60",
    x"60",x"60",x"77",x"00",x"B6",x"B6",x"B6",x"B6",x"B6",x"B6",x"B6",x"00",x"B6",x"00",x"60",x"60",
    x"60",x"60",x"77",x"00",x"77",x"B6",x"B6",x"00",x"B6",x"B6",x"B6",x"00",x"77",x"77",x"60",x"60",
    x"60",x"60",x"60",x"60",x"77",x"77",x"77",x"00",x"77",x"77",x"00",x"77",x"60",x"60",x"60",x"60",
    x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",

       --THE CRACKED ROCK OF GOLD
    x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",
    x"60",x"60",x"60",x"60",x"77",x"77",x"00",x"77",x"77",x"77",x"77",x"77",x"60",x"60",x"60",x"60",
    x"60",x"60",x"77",x"00",x"00",x"B6",x"00",x"B6",x"B6",x"B6",x"B6",x"00",x"77",x"77",x"60",x"60",
    x"60",x"60",x"77",x"B6",x"B6",x"00",x"00",x"B6",x"B6",x"00",x"00",x"B6",x"B6",x"77",x"60",x"60",
    x"60",x"77",x"00",x"B6",x"00",x"DD",x"B6",x"00",x"00",x"B6",x"B6",x"B6",x"B6",x"77",x"77",x"60",
    x"60",x"77",x"B6",x"00",x"B6",x"DD",x"B6",x"00",x"B6",x"DD",x"DD",x"B6",x"B6",x"00",x"00",x"60",
    x"60",x"77",x"B6",x"B6",x"DD",x"DD",x"00",x"B6",x"B6",x"B6",x"DD",x"DD",x"00",x"B6",x"77",x"60",
    x"60",x"77",x"B6",x"B6",x"DD",x"B6",x"00",x"B6",x"B6",x"B6",x"B6",x"00",x"00",x"B6",x"77",x"60",
    x"60",x"77",x"B6",x"B6",x"B6",x"B6",x"00",x"B6",x"B6",x"B6",x"B6",x"B6",x"DD",x"00",x"77",x"60",
    x"60",x"77",x"B6",x"B6",x"B6",x"00",x"DD",x"00",x"00",x"B6",x"B6",x"B6",x"B6",x"00",x"77",x"60",
    x"60",x"00",x"00",x"B6",x"B6",x"00",x"DD",x"B6",x"DD",x"00",x"DD",x"B6",x"00",x"B6",x"77",x"60",
    x"60",x"77",x"00",x"B6",x"00",x"B6",x"B6",x"B6",x"B6",x"B6",x"00",x"B6",x"00",x"77",x"77",x"60",
    x"60",x"60",x"77",x"00",x"B6",x"B6",x"B6",x"B6",x"B6",x"B6",x"B6",x"00",x"B6",x"00",x"60",x"60",
    x"60",x"60",x"77",x"00",x"77",x"B6",x"B6",x"00",x"B6",x"B6",x"B6",x"00",x"77",x"77",x"60",x"60",
    x"60",x"60",x"60",x"60",x"77",x"77",x"77",x"00",x"77",x"77",x"00",x"77",x"60",x"60",x"60",x"60",
    x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",

      --THE CRACKED ROCK OF greed
    x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",
    x"60",x"60",x"60",x"60",x"77",x"77",x"00",x"77",x"77",x"77",x"77",x"77",x"60",x"60",x"60",x"60",
    x"60",x"60",x"77",x"77",x"77",x"B6",x"00",x"B6",x"B6",x"B6",x"B6",x"00",x"77",x"77",x"60",x"60",
    x"60",x"60",x"00",x"00",x"B6",x"B6",x"00",x"B6",x"B6",x"00",x"00",x"B6",x"B6",x"77",x"60",x"60",
    x"60",x"77",x"77",x"B6",x"00",x"00",x"B6",x"00",x"00",x"E4",x"E4",x"B6",x"B6",x"77",x"77",x"60",
    x"60",x"00",x"B6",x"00",x"E4",x"B6",x"B6",x"00",x"E4",x"C0",x"C0",x"E4",x"B6",x"00",x"00",x"60",
    x"60",x"77",x"00",x"E4",x"C0",x"E4",x"00",x"B6",x"E4",x"C0",x"C0",x"E4",x"00",x"B6",x"77",x"60",
    x"60",x"77",x"B6",x"E4",x"C0",x"E4",x"00",x"B6",x"E4",x"C0",x"C0",x"00",x"00",x"B6",x"77",x"60",
    x"60",x"77",x"B6",x"B6",x"E4",x"B6",x"00",x"B6",x"B6",x"E4",x"E4",x"B6",x"B6",x"00",x"77",x"60",
    x"60",x"77",x"B6",x"B6",x"B6",x"00",x"B6",x"00",x"00",x"B6",x"B6",x"B6",x"B6",x"00",x"77",x"60",
    x"60",x"00",x"00",x"B6",x"B6",x"00",x"E4",x"E4",x"E4",x"00",x"B6",x"B6",x"00",x"B6",x"77",x"60",
    x"60",x"77",x"00",x"B6",x"00",x"E4",x"C0",x"C0",x"C0",x"E4",x"00",x"B6",x"00",x"7F",x"77",x"60",
    x"60",x"60",x"77",x"00",x"B6",x"B6",x"E4",x"E4",x"E4",x"B6",x"B6",x"00",x"B6",x"F7",x"60",x"60",
    x"60",x"60",x"77",x"00",x"77",x"B6",x"B6",x"00",x"B6",x"B6",x"B6",x"00",x"77",x"77",x"60",x"60",
    x"60",x"60",x"60",x"60",x"77",x"77",x"77",x"00",x"77",x"77",x"00",x"77",x"60",x"60",x"60",x"60",
    x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",x"60",



x"D0",x"D0",x"D0",x"D0",x"D1",x"D1",x"D1",x"D1",x"D2",x"D2",x"D2",x"D2",x"D3",x"D3",x"D3",x"D3",
x"D0",x"D0",x"D0",x"D0",x"D1",x"D1",x"D1",x"D1",x"D2",x"D2",x"D2",x"D2",x"D3",x"D3",x"D3",x"D3",
x"D0",x"D0",x"D0",x"D0",x"D1",x"D1",x"D1",x"D1",x"D2",x"D2",x"D2",x"D2",x"D3",x"D3",x"D3",x"D3",
x"D0",x"D0",x"D0",x"D0",x"D1",x"D1",x"D1",x"D1",x"D2",x"D2",x"D2",x"D2",x"D3",x"D3",x"D3",x"D3",
x"D4",x"D4",x"D4",x"D4",x"D5",x"D5",x"D5",x"D5",x"D6",x"D6",x"D6",x"D6",x"D7",x"D7",x"D7",x"D7",
x"D4",x"D4",x"D4",x"D4",x"D5",x"D5",x"D5",x"D5",x"D6",x"D6",x"D6",x"D6",x"D7",x"D7",x"D7",x"D7",
x"D4",x"D4",x"D4",x"D4",x"D5",x"D5",x"D5",x"D5",x"D6",x"D6",x"D6",x"D6",x"D7",x"D7",x"D7",x"D7",
x"D4",x"D4",x"D4",x"D4",x"D5",x"D5",x"D5",x"D5",x"D6",x"D6",x"D6",x"D6",x"D7",x"D7",x"D7",x"D7",
x"D8",x"D8",x"D8",x"D8",x"D9",x"D9",x"D9",x"D9",x"DA",x"DA",x"DA",x"DA",x"DB",x"DB",x"DB",x"DB",
x"D8",x"D8",x"D8",x"D8",x"D9",x"D9",x"D9",x"D9",x"DA",x"DA",x"DA",x"DA",x"DB",x"DB",x"DB",x"DB",
x"D8",x"D8",x"D8",x"D8",x"D9",x"D9",x"D9",x"D9",x"DA",x"DA",x"DA",x"DA",x"DB",x"DB",x"DB",x"DB",
x"D8",x"D8",x"D8",x"D8",x"D9",x"D9",x"D9",x"D9",x"DA",x"DA",x"DA",x"DA",x"DB",x"DB",x"DB",x"DB",
x"DC",x"DC",x"DC",x"DC",x"DD",x"DD",x"DD",x"DD",x"DE",x"DE",x"DE",x"DE",x"DF",x"DF",x"DF",x"DF",
x"DC",x"DC",x"DC",x"DC",x"DD",x"DD",x"DD",x"DD",x"DE",x"DE",x"DE",x"DE",x"DF",x"DF",x"DF",x"DF",
x"DC",x"DC",x"DC",x"DC",x"DD",x"DD",x"DD",x"DD",x"DE",x"DE",x"DE",x"DE",x"DF",x"DF",x"DF",x"DF",
x"DC",x"DC",x"DC",x"DC",x"DD",x"DD",x"DD",x"DD",x"DE",x"DE",x"DE",x"DE",x"DF",x"DF",x"DF",x"DF",


x"E0",x"E0",x"E0",x"E0",x"E1",x"E1",x"E1",x"E1",x"E2",x"E2",x"E2",x"E2",x"E3",x"E3",x"E3",x"E3",
x"E0",x"E0",x"E0",x"E0",x"E1",x"E1",x"E1",x"E1",x"E2",x"E2",x"E2",x"E2",x"E3",x"E3",x"E3",x"E3",
x"E0",x"E0",x"E0",x"E0",x"E1",x"E1",x"E1",x"E1",x"E2",x"E2",x"E2",x"E2",x"E3",x"E3",x"E3",x"E3",
x"E0",x"E0",x"E0",x"E0",x"E1",x"E1",x"E1",x"E1",x"E2",x"E2",x"E2",x"E2",x"E3",x"E3",x"E3",x"E3",
x"E4",x"E4",x"E4",x"E4",x"E5",x"E5",x"E5",x"E5",x"E6",x"E6",x"E6",x"E6",x"E7",x"E7",x"E7",x"E7",
x"E4",x"E4",x"E4",x"E4",x"E5",x"E5",x"E5",x"E5",x"E6",x"E6",x"E6",x"E6",x"E7",x"E7",x"E7",x"E7",
x"E4",x"E4",x"E4",x"E4",x"E5",x"E5",x"E5",x"E5",x"E6",x"E6",x"E6",x"E6",x"E7",x"E7",x"E7",x"E7",
x"E4",x"E4",x"E4",x"E4",x"E5",x"E5",x"E5",x"E5",x"E6",x"E6",x"E6",x"E6",x"E7",x"E7",x"E7",x"E7",
x"E8",x"E8",x"E8",x"E8",x"E9",x"E9",x"E9",x"E9",x"EA",x"EA",x"EA",x"EA",x"EB",x"EB",x"EB",x"EB",
x"E8",x"E8",x"E8",x"E8",x"E9",x"E9",x"E9",x"E9",x"EA",x"EA",x"EA",x"EA",x"EB",x"EB",x"EB",x"EB",
x"E8",x"E8",x"E8",x"E8",x"E9",x"E9",x"E9",x"E9",x"EA",x"EA",x"EA",x"EA",x"EB",x"EB",x"EB",x"EB",
x"E8",x"E8",x"E8",x"E8",x"E9",x"E9",x"E9",x"E9",x"EA",x"EA",x"EA",x"EA",x"EB",x"EB",x"EB",x"EB",
x"EC",x"EC",x"EC",x"EC",x"ED",x"ED",x"ED",x"ED",x"EE",x"EE",x"EE",x"EE",x"EF",x"EF",x"EF",x"EF",
x"EC",x"EC",x"EC",x"EC",x"ED",x"ED",x"ED",x"ED",x"EE",x"EE",x"EE",x"EE",x"EF",x"EF",x"EF",x"EF",
x"EC",x"EC",x"EC",x"EC",x"ED",x"ED",x"ED",x"ED",x"EE",x"EE",x"EE",x"EE",x"EF",x"EF",x"EF",x"EF",
x"EC",x"EC",x"EC",x"EC",x"ED",x"ED",x"ED",x"ED",x"EE",x"EE",x"EE",x"EE",x"EF",x"EF",x"EF",x"EF",


x"F0",x"F0",x"F0",x"F0",x"F1",x"F1",x"F1",x"F1",x"F2",x"F2",x"F2",x"F2",x"F3",x"F3",x"F3",x"F3",
x"F0",x"F0",x"F0",x"F0",x"F1",x"F1",x"F1",x"F1",x"F2",x"F2",x"F2",x"F2",x"F3",x"F3",x"F3",x"F3",
x"F0",x"F0",x"F0",x"F0",x"F1",x"F1",x"F1",x"F1",x"F2",x"F2",x"F2",x"F2",x"F3",x"F3",x"F3",x"F3",
x"F0",x"F0",x"F0",x"F0",x"F1",x"F1",x"F1",x"F1",x"F2",x"F2",x"F2",x"F2",x"F3",x"F3",x"F3",x"F3",
x"F4",x"F4",x"F4",x"F4",x"F5",x"F5",x"F5",x"F5",x"F6",x"F6",x"F6",x"F6",x"F7",x"F7",x"F7",x"F7",
x"F4",x"F4",x"F4",x"F4",x"F5",x"F5",x"F5",x"F5",x"F6",x"F6",x"F6",x"F6",x"F7",x"F7",x"F7",x"F7",
x"F4",x"F4",x"F4",x"F4",x"F5",x"F5",x"F5",x"F5",x"F6",x"F6",x"F6",x"F6",x"F7",x"F7",x"F7",x"F7",
x"F4",x"F4",x"F4",x"F4",x"F5",x"F5",x"F5",x"F5",x"F6",x"F6",x"F6",x"F6",x"F7",x"F7",x"F7",x"F7",
x"F8",x"F8",x"F8",x"F8",x"F9",x"F9",x"F9",x"F9",x"FA",x"FA",x"FA",x"FA",x"FB",x"FB",x"FB",x"FB",
x"F8",x"F8",x"F8",x"F8",x"F9",x"F9",x"F9",x"F9",x"FA",x"FA",x"FA",x"FA",x"FB",x"FB",x"FB",x"FB",
x"F8",x"F8",x"F8",x"F8",x"F9",x"F9",x"F9",x"F9",x"FA",x"FA",x"FA",x"FA",x"FB",x"FB",x"FB",x"FB",
x"F8",x"F8",x"F8",x"F8",x"F9",x"F9",x"F9",x"F9",x"FA",x"FA",x"FA",x"FA",x"FB",x"FB",x"FB",x"FB",
x"FC",x"FC",x"FC",x"FC",x"FD",x"FD",x"FD",x"FD",x"FE",x"FE",x"FE",x"FE",x"FF",x"FF",x"FF",x"FF",
x"FC",x"FC",x"FC",x"FC",x"FD",x"FD",x"FD",x"FD",x"FE",x"FE",x"FE",x"FE",x"FF",x"FF",x"FF",x"FF",
x"FC",x"FC",x"FC",x"FC",x"FD",x"FD",x"FD",x"FD",x"FE",x"FE",x"FE",x"FE",x"FF",x"FF",x"FF",x"FF",
x"FC",x"FC",x"FC",x"FC",x"FD",x"FD",x"FD",x"FD",x"FE",x"FE",x"FE",x"FE",x"FF",x"FF",x"FF",x"FF",


    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
   
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",     

    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",

    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",

    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",


    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",

    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",

    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",

    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",

    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",

    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",

    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",

    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",

    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",

    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",

    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",

    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",

    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",

    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",

    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",

    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",

    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",

    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",

    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",

    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",

    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",

    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
    x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",

    x"00",x"10",x"20",x"30",x"40",x"50",x"60",x"70",x"80",x"90",x"A0",x"B0",x"C0",x"D0",x"E0",x"F0", 
    x"00",x"11",x"21",x"31",x"41",x"51",x"61",x"71",x"81",x"91",x"A1",x"B1",x"C1",x"D1",x"E1",x"F1",
    x"00",x"12",x"22",x"32",x"42",x"52",x"62",x"72",x"82",x"92",x"A2",x"B2",x"C2",x"D2",x"E2",x"F2",
    x"00",x"13",x"23",x"33",x"77",x"53",x"63",x"DF",x"83",x"93",x"A3",x"B3",x"C3",x"D3",x"E3",x"F3",
    x"04",x"14",x"24",x"34",x"44",x"54",x"64",x"74",x"84",x"94",x"A4",x"B4",x"C4",x"D4",x"E4",x"F4",
    x"05",x"15",x"25",x"35",x"45",x"55",x"65",x"75",x"85",x"95",x"A5",x"B5",x"C5",x"D5",x"E5",x"F5",
    x"06",x"16",x"26",x"36",x"46",x"56",x"66",x"76",x"86",x"96",x"A6",x"B6",x"C6",x"D6",x"E6",x"F6",
    x"07",x"17",x"27",x"37",x"47",x"57",x"67",x"DF",x"87",x"97",x"A7",x"B7",x"C7",x"D7",x"E7",x"F7",
    x"08",x"18",x"28",x"38",x"48",x"58",x"68",x"78",x"88",x"98",x"A8",x"B8",x"C8",x"D8",x"E8",x"F8",
    x"09",x"19",x"29",x"39",x"49",x"59",x"69",x"79",x"89",x"99",x"A9",x"B9",x"C9",x"D9",x"E9",x"F9",
    x"0A",x"1A",x"2A",x"3A",x"4A",x"5A",x"6A",x"7A",x"8A",x"9A",x"AA",x"BA",x"CA",x"DA",x"EA",x"FA",
    x"0B",x"1B",x"2B",x"3B",x"4B",x"5B",x"6B",x"7B",x"8B",x"9B",x"AB",x"BB",x"CB",x"DB",x"EB",x"FB",
    x"0C",x"1C",x"2C",x"3C",x"4C",x"5C",x"6C",x"7C",x"8C",x"9C",x"AC",x"BC",x"CC",x"DC",x"EC",x"FC",
    x"0D",x"1D",x"2D",x"3D",x"4D",x"5D",x"6D",x"7D",x"8D",x"9D",x"AD",x"BD",x"CD",x"DD",x"ED",x"FD",
    x"0E",x"1E",x"2E",x"3E",x"4E",x"5E",x"6E",x"7E",x"8E",x"9E",x"AE",x"BE",x"CE",x"DE",x"EE",x"FE",
    x"0F",x"1F",x"2F",x"3F",x"4F",x"5F",x"6F",x"7F",x"8F",x"9F",x"AF",x"BF",x"CF",x"DF",x"EF",x"FF"
    );

begin
    pixel_out <= tMem( (to_integer(tile_index) * 256) + (to_integer(tile_pixel_Y) * 16) + to_integer(tile_pixel_X) );
end Behavioral;
